`timescale 1ns / 1ps
// Copyright 2017 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the “License�?); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an “AS IS�? BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );


//   const logic [0:472] [31:0] mem = {

// 32'h44054101,
// 32'h91220436,
// 32'h04524405,
// 32'h44019122,
// 32'hCE86711D,
// 32'h1080CCA2,
// 32'h29954505,
// 32'h04000593,
// 32'h2E894501,
// 32'hFE042623,
// 32'h0001A039,
// 32'hFEC42783,
// 32'h26230785,
// 32'h2703FEF4,
// 32'h6785FEC4,
// 32'hBB778793,
// 32'hFEE7D5E3,
// 32'h1A1027B7,
// 32'h07130791,
// 32'hC3980200,
// 32'h87AA2A5D,
// 32'h0593CB81,
// 32'h67C10240,
// 32'h6CC78513,
// 32'hA0012645,
// 32'h67C145C5,
// 32'h6F478513,
// 32'h24232E51,
// 32'h4581FE04,
// 32'h29D54501,
// 32'hFE842783,
// 32'h069307A2,
// 32'h863E0200,
// 32'h454D45A1,
// 32'h0513298D,
// 32'h2B011000,
// 32'h45014581,
// 32'h079323B9,
// 32'h0593FA04,
// 32'h853E1000,
// 32'h27832345,
// 32'h2A23FA04,
// 32'h2783FCF4,
// 32'h2223FA44,
// 32'h2783FEF4,
// 32'h2823FA84,
// 32'h2783FCF4,
// 32'h2623FAC4,
// 32'h2783FCF4,
// 32'h2423FB04,
// 32'h2783FCF4,
// 32'h2023FB44,
// 32'h2783FEF4,
// 32'h2223FB84,
// 32'h2783FCF4,
// 32'h2023FBC4,
// 32'h45D5FCF4,
// 32'h851367C1,
// 32'h2E197087,
// 32'hFD442783,
// 32'hFEF42423,
// 32'hFC042E23,
// 32'h2783A881,
// 32'h07A2FE84,
// 32'h02000693,
// 32'h45A1863E,
// 32'h2EC5454D,
// 32'h29416521,
// 32'h45014581,
// 32'h65A121F9,
// 32'hFE442503,
// 32'h27032315,
// 32'h6785FE44,
// 32'h222397BA,
// 32'h2703FEF4,
// 32'h6785FE84,
// 32'h242397BA,
// 32'h2783FEF4,
// 32'h853EFDC4,
// 32'h27832AB5,
// 32'h0785FDC4,
// 32'hFCF42E23,
// 32'hFDC42703,
// 32'hFCC42783,
// 32'hFAF745E3,
// 32'h21F90001,
// 32'h67C1872A,
// 32'h8F7D17FD,
// 32'h1AE34785,
// 32'h45B5FEF7,
// 32'h851367C1,
// 32'h2C497207,
// 32'h27832601,
// 32'h2423FC84,
// 32'h2C23FEF4,
// 32'hA889FC04,
// 32'hFE842783,
// 32'h069307A2,
// 32'h863E0200,
// 32'h051345A1,
// 32'h26A50EB0,
// 32'h21216521,
// 32'h45094581,
// 32'h65A12199,
// 32'hFE042503,
// 32'h27032971,
// 32'h6785FE04,
// 32'h202397BA,
// 32'h2703FEF4,
// 32'h6785FE84,
// 32'h242397BA,
// 32'h2783FEF4,
// 32'h853EFD84,
// 32'h278328D5,
// 32'h0785FD84,
// 32'hFCF42C23,
// 32'hFD842703,
// 32'hFC042783,
// 32'hFAF744E3,
// 32'h02200593,
// 32'h851367C1,
// 32'h2C297307,
// 32'h77B72461,
// 32'h07A11A10,
// 32'h0007A023,
// 32'h08000513,
// 32'h47812045,
// 32'h40F6853E,
// 32'h61254466,
// 32'h11018082,
// 32'hCC22CE06,
// 32'h26231000,
// 32'h4681FE04,
// 32'h45A14601,
// 32'h09F00513,
// 32'h05132CF9,
// 32'h2EB50400,
// 32'h45014581,
// 32'h45812689,
// 32'h2E554501,
// 32'hFE440793,
// 32'h04000593,
// 32'h2119853E,
// 32'hFE442783,
// 32'h0187D713,
// 32'h07634785,
// 32'h278300F7,
// 32'h0785FEC4,
// 32'hFEF42623,
// 32'hFE442783,
// 32'h4087D713,
// 32'h17FD67C1,
// 32'h07938F7D,
// 32'h02632190,
// 32'h278302F7,
// 32'hD713FE44,
// 32'h67C14087,
// 32'h8F7D17FD,
// 32'h07E16789,
// 32'h00F70763,
// 32'hFEC42783,
// 32'h26230785,
// 32'h2783FEF4,
// 32'h853EFEC4,
// 32'h446240F2,
// 32'h80826105,
// 32'hCE221101,
// 32'h26231000,
// 32'h2783FEA4,
// 32'h8067FEC4,
// 32'h00010007,
// 32'h00010001,
// 32'h44720001,
// 32'h80826105,
// 32'hD6067179,
// 32'h1800D422,
// 32'hFCA42E23,
// 32'hFDC42783,
// 32'h26238BBD,
// 32'h2783FEF4,
// 32'h8391FDC4,
// 32'hFEF42423,
// 32'h67C14599,
// 32'h75478513,
// 32'h27032205,
// 32'h67C1FE84,
// 32'h6BC78793,
// 32'h458597BA,
// 32'h2239853E,
// 32'hFEC42703,
// 32'h879367C1,
// 32'h97BA6BC7,
// 32'h853E4585,
// 32'h459928F5,
// 32'h851367C1,
// 32'h28CD75C7,
// 32'h00012285,
// 32'h542250B2,
// 32'h80826145,
// 32'hD6227179,
// 32'h2E231800,
// 32'h2C23FCA4,
// 32'h77B7FCB4,
// 32'h439C1A10,
// 32'hFEF42623,
// 32'h27834705,
// 32'h17B3FDC4,
// 32'hC71300F7,
// 32'h2783FFF7,
// 32'h8FF9FEC4,
// 32'hFEF42623,
// 32'hFD842703,
// 32'hFDC42783,
// 32'h00F71733,
// 32'hFEC42783,
// 32'h26238FD9,
// 32'h77B7FEF4,
// 32'h27031A10,
// 32'hC398FEC4,
// 32'h54320001,
// 32'h80826145,
// 32'hCE221101,
// 32'h26231000,
// 32'h87AEFEA4,
// 32'hFEF41523,
// 32'h1A1077B7,
// 32'h43980791,
// 32'h1A1077B7,
// 32'h67130791,
// 32'hC3980027,
// 32'h1A1007B7,
// 32'h071307B1,
// 32'hC3980830,
// 32'hFEA45783,
// 32'h07C283A1,
// 32'h873E83C1,
// 32'h1A1007B7,
// 32'h77130791,
// 32'hC3980FF7,
// 32'hFEA45703,
// 32'h1A1007B7,
// 32'h0FF77713,
// 32'h07B7C398,
// 32'h07A11A10,
// 32'h0A700713,
// 32'h07B7C398,
// 32'h07B11A10,
// 32'hC398470D,
// 32'h1A1007B7,
// 32'h439C0791,
// 32'h0F07F713,
// 32'h1A1007B7,
// 32'h67130791,
// 32'hC3980027,
// 32'h44720001,
// 32'h80826105,
// 32'hD6227179,
// 32'h2E231800,
// 32'h2C23FCA4,
// 32'hA891FCB4,
// 32'h07B70001,
// 32'h07D11A10,
// 32'hF793439C,
// 32'hDBF50207,
// 32'hFE042623,
// 32'h2783A035,
// 32'h8713FDC4,
// 32'h2E230017,
// 32'hC703FCE4,
// 32'h07B70007,
// 32'hC3981A10,
// 32'hFD842783,
// 32'h2C2317FD,
// 32'h2783FCF4,
// 32'h0785FEC4,
// 32'hFEF42623,
// 32'hFEC42703,
// 32'h03F00793,
// 32'h00E7E563,
// 32'hFD842783,
// 32'h2783F3F9,
// 32'hF7CDFD84,
// 32'h54320001,
// 32'h80826145,
// 32'hC6221141,
// 32'h00010800,
// 32'h1A1007B7,
// 32'h439C07D1,
// 32'h0407F793,
// 32'h0001DBF5,
// 32'h01414432,
// 32'h11018082,
// 32'hCC22CE06,
// 32'h26231000,
// 32'h4581FEA4,
// 32'h3DBD453D,
// 32'h45394581,
// 32'h45813DA5,
// 32'h3D8D4535,
// 32'h45314581,
// 32'h278335B5,
// 32'h5563FEC4,
// 32'h458100F0,
// 32'h3DB94541,
// 32'hFEC42703,
// 32'hD5634785,
// 32'h458100E7,
// 32'h35B9452D,
// 32'hFEC42703,
// 32'hD5634789,
// 32'h458100E7,
// 32'h3D3D4501,
// 32'hFEC42703,
// 32'hD563478D,
// 32'h458100E7,
// 32'h353D4505,
// 32'h40F20001,
// 32'h61054462,
// 32'h71798082,
// 32'h1800D622,
// 32'hFCA42E23,
// 32'hFCB42C23,
// 32'hFCC42A23,
// 32'hFCD42823,
// 32'h02000713,
// 32'hFD842783,
// 32'h40F707B3,
// 32'hFDC42703,
// 32'h00F717B3,
// 32'hFEF42623,
// 32'h1A1027B7,
// 32'h270307A1,
// 32'hC398FEC4,
// 32'h1A1027B7,
// 32'h270307B1,
// 32'hC398FD44,
// 32'hFD842783,
// 32'h03F7F693,
// 32'hFD042783,
// 32'h00879713,
// 32'h87936791,
// 32'h8F7DF007,
// 32'h1A1027B7,
// 32'h8F5507C1,
// 32'h0001C398,
// 32'h61455432,
// 32'h11018082,
// 32'h1000CE22,
// 32'hFEA42623,
// 32'hFEB42423,
// 32'hFE842783,
// 32'h86BE07C2,
// 32'hFEC42703,
// 32'h17FD67C1,
// 32'hE7338FF9,
// 32'h27B700F6,
// 32'h07D11A10,
// 32'h0001C398,
// 32'h61054472,
// 32'h71798082,
// 32'h1800D622,
// 32'hFCA42E23,
// 32'h1A1027B7,
// 32'h439C07C1,
// 32'hFEF42623,
// 32'hFDC42783,
// 32'h873E07C2,
// 32'hFEC42783,
// 32'h67C186BE,
// 32'h8FF517FD,
// 32'h26238FD9,
// 32'h27B7FEF4,
// 32'h07C11A10,
// 32'hFEC42703,
// 32'h0001C398,
// 32'h61455432,
// 32'h11018082,
// 32'h1000CE22,
// 32'hFEA42623,
// 32'hFEB42423,
// 32'hFE842783,
// 32'h470507A1,
// 32'h00F71733,
// 32'h87936785,
// 32'h76B3F007,
// 32'h470500F7,
// 32'hFEC42783,
// 32'h00F717B3,
// 32'h0FF7F713,
// 32'h1A1027B7,
// 32'hC3988F55,
// 32'h44720001,
// 32'h80826105,
// 32'hCE221101,
// 32'h27B71000,
// 32'h439C1A10,
// 32'hFEF42623,
// 32'hFEC42783,
// 32'h4472853E,
// 32'h80826105,
// 32'hD6227179,
// 32'h2E231800,
// 32'h2C23FCA4,
// 32'h2783FCB4,
// 32'h8795FD84,
// 32'h7FF7F793,
// 32'hFEF42623,
// 32'hFD842783,
// 32'hC7918BFD,
// 32'hFEC42783,
// 32'h26230785,
// 32'h2423FEF4,
// 32'hA815FE04,
// 32'h27B70001,
// 32'h439C1A10,
// 32'hF79387C1,
// 32'hDBF50FF7,
// 32'h1A1027B7,
// 32'h02078713,
// 32'hFE842783,
// 32'h2683078A,
// 32'h97B6FDC4,
// 32'hC3984318,
// 32'hFE842783,
// 32'h24230785,
// 32'h2703FEF4,
// 32'h2783FE84,
// 32'h43E3FEC4,
// 32'h0001FCF7,
// 32'h61455432,
// 32'h31308082,
// 32'h35343332,
// 32'h39383736,
// 32'h44434241,
// 32'h52454645,
// 32'h3A524F52,
// 32'h61705320,
// 32'h6F69736E,
// 32'h5053206E,
// 32'h6C662049,
// 32'h20687361,
// 32'h20746F6E,
// 32'h6E756F66,
// 32'h00000A64,
// 32'h6F4C0000,
// 32'h6E696461,
// 32'h72662067,
// 32'h53206D6F,
// 32'h000A4950,
// 32'h6F430000,
// 32'h6E697970,
// 32'h6E492067,
// 32'h75727473,
// 32'h6F697463,
// 32'h000A736E,
// 32'h6F430000,
// 32'h6E697970,
// 32'h61442067,
// 32'h000A6174,
// 32'h6F440000,
// 32'h202C656E,
// 32'h706D756A,
// 32'h20676E69,
// 32'h49206F74,
// 32'h7274736E,
// 32'h69746375,
// 32'h52206E6F,
// 32'h0A2E4D41,
// 32'h6C420000,
// 32'h206B636F,
// 32'h64200000,
// 32'h0A656E6F,
// 32'h0000C600

//     };

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end


  // assign Q = mem[A_Q];


endmodule