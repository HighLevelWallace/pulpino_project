
module decoder_8to256(
	input  [  7:0] addr_i,
	output [255:0] select_o
);

assign select_o[0] = (addr_i == 8'd0) ? 1 : 0;
assign select_o[1] = (addr_i == 8'd1) ? 1 : 0;
assign select_o[2] = (addr_i == 8'd2) ? 1 : 0;
assign select_o[3] = (addr_i == 8'd3) ? 1 : 0;
assign select_o[4] = (addr_i == 8'd4) ? 1 : 0;
assign select_o[5] = (addr_i == 8'd5) ? 1 : 0;
assign select_o[6] = (addr_i == 8'd6) ? 1 : 0;
assign select_o[7] = (addr_i == 8'd7) ? 1 : 0;
assign select_o[8] = (addr_i == 8'd8) ? 1 : 0;
assign select_o[9] = (addr_i == 8'd9) ? 1 : 0;
assign select_o[10] = (addr_i == 8'd10) ? 1 : 0;
assign select_o[11] = (addr_i == 8'd11) ? 1 : 0;
assign select_o[12] = (addr_i == 8'd12) ? 1 : 0;
assign select_o[13] = (addr_i == 8'd13) ? 1 : 0;
assign select_o[14] = (addr_i == 8'd14) ? 1 : 0;
assign select_o[15] = (addr_i == 8'd15) ? 1 : 0;
assign select_o[16] = (addr_i == 8'd16) ? 1 : 0;
assign select_o[17] = (addr_i == 8'd17) ? 1 : 0;
assign select_o[18] = (addr_i == 8'd18) ? 1 : 0;
assign select_o[19] = (addr_i == 8'd19) ? 1 : 0;
assign select_o[20] = (addr_i == 8'd20) ? 1 : 0;
assign select_o[21] = (addr_i == 8'd21) ? 1 : 0;
assign select_o[22] = (addr_i == 8'd22) ? 1 : 0;
assign select_o[23] = (addr_i == 8'd23) ? 1 : 0;
assign select_o[24] = (addr_i == 8'd24) ? 1 : 0;
assign select_o[25] = (addr_i == 8'd25) ? 1 : 0;
assign select_o[26] = (addr_i == 8'd26) ? 1 : 0;
assign select_o[27] = (addr_i == 8'd27) ? 1 : 0;
assign select_o[28] = (addr_i == 8'd28) ? 1 : 0;
assign select_o[29] = (addr_i == 8'd29) ? 1 : 0;
assign select_o[30] = (addr_i == 8'd30) ? 1 : 0;
assign select_o[31] = (addr_i == 8'd31) ? 1 : 0;
assign select_o[32] = (addr_i == 8'd32) ? 1 : 0;
assign select_o[33] = (addr_i == 8'd33) ? 1 : 0;
assign select_o[34] = (addr_i == 8'd34) ? 1 : 0;
assign select_o[35] = (addr_i == 8'd35) ? 1 : 0;
assign select_o[36] = (addr_i == 8'd36) ? 1 : 0;
assign select_o[37] = (addr_i == 8'd37) ? 1 : 0;
assign select_o[38] = (addr_i == 8'd38) ? 1 : 0;
assign select_o[39] = (addr_i == 8'd39) ? 1 : 0;
assign select_o[40] = (addr_i == 8'd40) ? 1 : 0;
assign select_o[41] = (addr_i == 8'd41) ? 1 : 0;
assign select_o[42] = (addr_i == 8'd42) ? 1 : 0;
assign select_o[43] = (addr_i == 8'd43) ? 1 : 0;
assign select_o[44] = (addr_i == 8'd44) ? 1 : 0;
assign select_o[45] = (addr_i == 8'd45) ? 1 : 0;
assign select_o[46] = (addr_i == 8'd46) ? 1 : 0;
assign select_o[47] = (addr_i == 8'd47) ? 1 : 0;
assign select_o[48] = (addr_i == 8'd48) ? 1 : 0;
assign select_o[49] = (addr_i == 8'd49) ? 1 : 0;
assign select_o[50] = (addr_i == 8'd50) ? 1 : 0;
assign select_o[51] = (addr_i == 8'd51) ? 1 : 0;
assign select_o[52] = (addr_i == 8'd52) ? 1 : 0;
assign select_o[53] = (addr_i == 8'd53) ? 1 : 0;
assign select_o[54] = (addr_i == 8'd54) ? 1 : 0;
assign select_o[55] = (addr_i == 8'd55) ? 1 : 0;
assign select_o[56] = (addr_i == 8'd56) ? 1 : 0;
assign select_o[57] = (addr_i == 8'd57) ? 1 : 0;
assign select_o[58] = (addr_i == 8'd58) ? 1 : 0;
assign select_o[59] = (addr_i == 8'd59) ? 1 : 0;
assign select_o[60] = (addr_i == 8'd60) ? 1 : 0;
assign select_o[61] = (addr_i == 8'd61) ? 1 : 0;
assign select_o[62] = (addr_i == 8'd62) ? 1 : 0;
assign select_o[63] = (addr_i == 8'd63) ? 1 : 0;
assign select_o[64] = (addr_i == 8'd64) ? 1 : 0;
assign select_o[65] = (addr_i == 8'd65) ? 1 : 0;
assign select_o[66] = (addr_i == 8'd66) ? 1 : 0;
assign select_o[67] = (addr_i == 8'd67) ? 1 : 0;
assign select_o[68] = (addr_i == 8'd68) ? 1 : 0;
assign select_o[69] = (addr_i == 8'd69) ? 1 : 0;
assign select_o[70] = (addr_i == 8'd70) ? 1 : 0;
assign select_o[71] = (addr_i == 8'd71) ? 1 : 0;
assign select_o[72] = (addr_i == 8'd72) ? 1 : 0;
assign select_o[73] = (addr_i == 8'd73) ? 1 : 0;
assign select_o[74] = (addr_i == 8'd74) ? 1 : 0;
assign select_o[75] = (addr_i == 8'd75) ? 1 : 0;
assign select_o[76] = (addr_i == 8'd76) ? 1 : 0;
assign select_o[77] = (addr_i == 8'd77) ? 1 : 0;
assign select_o[78] = (addr_i == 8'd78) ? 1 : 0;
assign select_o[79] = (addr_i == 8'd79) ? 1 : 0;
assign select_o[80] = (addr_i == 8'd80) ? 1 : 0;
assign select_o[81] = (addr_i == 8'd81) ? 1 : 0;
assign select_o[82] = (addr_i == 8'd82) ? 1 : 0;
assign select_o[83] = (addr_i == 8'd83) ? 1 : 0;
assign select_o[84] = (addr_i == 8'd84) ? 1 : 0;
assign select_o[85] = (addr_i == 8'd85) ? 1 : 0;
assign select_o[86] = (addr_i == 8'd86) ? 1 : 0;
assign select_o[87] = (addr_i == 8'd87) ? 1 : 0;
assign select_o[88] = (addr_i == 8'd88) ? 1 : 0;
assign select_o[89] = (addr_i == 8'd89) ? 1 : 0;
assign select_o[90] = (addr_i == 8'd90) ? 1 : 0;
assign select_o[91] = (addr_i == 8'd91) ? 1 : 0;
assign select_o[92] = (addr_i == 8'd92) ? 1 : 0;
assign select_o[93] = (addr_i == 8'd93) ? 1 : 0;
assign select_o[94] = (addr_i == 8'd94) ? 1 : 0;
assign select_o[95] = (addr_i == 8'd95) ? 1 : 0;
assign select_o[96] = (addr_i == 8'd96) ? 1 : 0;
assign select_o[97] = (addr_i == 8'd97) ? 1 : 0;
assign select_o[98] = (addr_i == 8'd98) ? 1 : 0;
assign select_o[99] = (addr_i == 8'd99) ? 1 : 0;
assign select_o[100] = (addr_i == 8'd100) ? 1 : 0;
assign select_o[101] = (addr_i == 8'd101) ? 1 : 0;
assign select_o[102] = (addr_i == 8'd102) ? 1 : 0;
assign select_o[103] = (addr_i == 8'd103) ? 1 : 0;
assign select_o[104] = (addr_i == 8'd104) ? 1 : 0;
assign select_o[105] = (addr_i == 8'd105) ? 1 : 0;
assign select_o[106] = (addr_i == 8'd106) ? 1 : 0;
assign select_o[107] = (addr_i == 8'd107) ? 1 : 0;
assign select_o[108] = (addr_i == 8'd108) ? 1 : 0;
assign select_o[109] = (addr_i == 8'd109) ? 1 : 0;
assign select_o[110] = (addr_i == 8'd110) ? 1 : 0;
assign select_o[111] = (addr_i == 8'd111) ? 1 : 0;
assign select_o[112] = (addr_i == 8'd112) ? 1 : 0;
assign select_o[113] = (addr_i == 8'd113) ? 1 : 0;
assign select_o[114] = (addr_i == 8'd114) ? 1 : 0;
assign select_o[115] = (addr_i == 8'd115) ? 1 : 0;
assign select_o[116] = (addr_i == 8'd116) ? 1 : 0;
assign select_o[117] = (addr_i == 8'd117) ? 1 : 0;
assign select_o[118] = (addr_i == 8'd118) ? 1 : 0;
assign select_o[119] = (addr_i == 8'd119) ? 1 : 0;
assign select_o[120] = (addr_i == 8'd120) ? 1 : 0;
assign select_o[121] = (addr_i == 8'd121) ? 1 : 0;
assign select_o[122] = (addr_i == 8'd122) ? 1 : 0;
assign select_o[123] = (addr_i == 8'd123) ? 1 : 0;
assign select_o[124] = (addr_i == 8'd124) ? 1 : 0;
assign select_o[125] = (addr_i == 8'd125) ? 1 : 0;
assign select_o[126] = (addr_i == 8'd126) ? 1 : 0;
assign select_o[127] = (addr_i == 8'd127) ? 1 : 0;
assign select_o[128] = (addr_i == 8'd128) ? 1 : 0;
assign select_o[129] = (addr_i == 8'd129) ? 1 : 0;
assign select_o[130] = (addr_i == 8'd130) ? 1 : 0;
assign select_o[131] = (addr_i == 8'd131) ? 1 : 0;
assign select_o[132] = (addr_i == 8'd132) ? 1 : 0;
assign select_o[133] = (addr_i == 8'd133) ? 1 : 0;
assign select_o[134] = (addr_i == 8'd134) ? 1 : 0;
assign select_o[135] = (addr_i == 8'd135) ? 1 : 0;
assign select_o[136] = (addr_i == 8'd136) ? 1 : 0;
assign select_o[137] = (addr_i == 8'd137) ? 1 : 0;
assign select_o[138] = (addr_i == 8'd138) ? 1 : 0;
assign select_o[139] = (addr_i == 8'd139) ? 1 : 0;
assign select_o[140] = (addr_i == 8'd140) ? 1 : 0;
assign select_o[141] = (addr_i == 8'd141) ? 1 : 0;
assign select_o[142] = (addr_i == 8'd142) ? 1 : 0;
assign select_o[143] = (addr_i == 8'd143) ? 1 : 0;
assign select_o[144] = (addr_i == 8'd144) ? 1 : 0;
assign select_o[145] = (addr_i == 8'd145) ? 1 : 0;
assign select_o[146] = (addr_i == 8'd146) ? 1 : 0;
assign select_o[147] = (addr_i == 8'd147) ? 1 : 0;
assign select_o[148] = (addr_i == 8'd148) ? 1 : 0;
assign select_o[149] = (addr_i == 8'd149) ? 1 : 0;
assign select_o[150] = (addr_i == 8'd150) ? 1 : 0;
assign select_o[151] = (addr_i == 8'd151) ? 1 : 0;
assign select_o[152] = (addr_i == 8'd152) ? 1 : 0;
assign select_o[153] = (addr_i == 8'd153) ? 1 : 0;
assign select_o[154] = (addr_i == 8'd154) ? 1 : 0;
assign select_o[155] = (addr_i == 8'd155) ? 1 : 0;
assign select_o[156] = (addr_i == 8'd156) ? 1 : 0;
assign select_o[157] = (addr_i == 8'd157) ? 1 : 0;
assign select_o[158] = (addr_i == 8'd158) ? 1 : 0;
assign select_o[159] = (addr_i == 8'd159) ? 1 : 0;
assign select_o[160] = (addr_i == 8'd160) ? 1 : 0;
assign select_o[161] = (addr_i == 8'd161) ? 1 : 0;
assign select_o[162] = (addr_i == 8'd162) ? 1 : 0;
assign select_o[163] = (addr_i == 8'd163) ? 1 : 0;
assign select_o[164] = (addr_i == 8'd164) ? 1 : 0;
assign select_o[165] = (addr_i == 8'd165) ? 1 : 0;
assign select_o[166] = (addr_i == 8'd166) ? 1 : 0;
assign select_o[167] = (addr_i == 8'd167) ? 1 : 0;
assign select_o[168] = (addr_i == 8'd168) ? 1 : 0;
assign select_o[169] = (addr_i == 8'd169) ? 1 : 0;
assign select_o[170] = (addr_i == 8'd170) ? 1 : 0;
assign select_o[171] = (addr_i == 8'd171) ? 1 : 0;
assign select_o[172] = (addr_i == 8'd172) ? 1 : 0;
assign select_o[173] = (addr_i == 8'd173) ? 1 : 0;
assign select_o[174] = (addr_i == 8'd174) ? 1 : 0;
assign select_o[175] = (addr_i == 8'd175) ? 1 : 0;
assign select_o[176] = (addr_i == 8'd176) ? 1 : 0;
assign select_o[177] = (addr_i == 8'd177) ? 1 : 0;
assign select_o[178] = (addr_i == 8'd178) ? 1 : 0;
assign select_o[179] = (addr_i == 8'd179) ? 1 : 0;
assign select_o[180] = (addr_i == 8'd180) ? 1 : 0;
assign select_o[181] = (addr_i == 8'd181) ? 1 : 0;
assign select_o[182] = (addr_i == 8'd182) ? 1 : 0;
assign select_o[183] = (addr_i == 8'd183) ? 1 : 0;
assign select_o[184] = (addr_i == 8'd184) ? 1 : 0;
assign select_o[185] = (addr_i == 8'd185) ? 1 : 0;
assign select_o[186] = (addr_i == 8'd186) ? 1 : 0;
assign select_o[187] = (addr_i == 8'd187) ? 1 : 0;
assign select_o[188] = (addr_i == 8'd188) ? 1 : 0;
assign select_o[189] = (addr_i == 8'd189) ? 1 : 0;
assign select_o[190] = (addr_i == 8'd190) ? 1 : 0;
assign select_o[191] = (addr_i == 8'd191) ? 1 : 0;
assign select_o[192] = (addr_i == 8'd192) ? 1 : 0;
assign select_o[193] = (addr_i == 8'd193) ? 1 : 0;
assign select_o[194] = (addr_i == 8'd194) ? 1 : 0;
assign select_o[195] = (addr_i == 8'd195) ? 1 : 0;
assign select_o[196] = (addr_i == 8'd196) ? 1 : 0;
assign select_o[197] = (addr_i == 8'd197) ? 1 : 0;
assign select_o[198] = (addr_i == 8'd198) ? 1 : 0;
assign select_o[199] = (addr_i == 8'd199) ? 1 : 0;
assign select_o[200] = (addr_i == 8'd200) ? 1 : 0;
assign select_o[201] = (addr_i == 8'd201) ? 1 : 0;
assign select_o[202] = (addr_i == 8'd202) ? 1 : 0;
assign select_o[203] = (addr_i == 8'd203) ? 1 : 0;
assign select_o[204] = (addr_i == 8'd204) ? 1 : 0;
assign select_o[205] = (addr_i == 8'd205) ? 1 : 0;
assign select_o[206] = (addr_i == 8'd206) ? 1 : 0;
assign select_o[207] = (addr_i == 8'd207) ? 1 : 0;
assign select_o[208] = (addr_i == 8'd208) ? 1 : 0;
assign select_o[209] = (addr_i == 8'd209) ? 1 : 0;
assign select_o[210] = (addr_i == 8'd210) ? 1 : 0;
assign select_o[211] = (addr_i == 8'd211) ? 1 : 0;
assign select_o[212] = (addr_i == 8'd212) ? 1 : 0;
assign select_o[213] = (addr_i == 8'd213) ? 1 : 0;
assign select_o[214] = (addr_i == 8'd214) ? 1 : 0;
assign select_o[215] = (addr_i == 8'd215) ? 1 : 0;
assign select_o[216] = (addr_i == 8'd216) ? 1 : 0;
assign select_o[217] = (addr_i == 8'd217) ? 1 : 0;
assign select_o[218] = (addr_i == 8'd218) ? 1 : 0;
assign select_o[219] = (addr_i == 8'd219) ? 1 : 0;
assign select_o[220] = (addr_i == 8'd220) ? 1 : 0;
assign select_o[221] = (addr_i == 8'd221) ? 1 : 0;
assign select_o[222] = (addr_i == 8'd222) ? 1 : 0;
assign select_o[223] = (addr_i == 8'd223) ? 1 : 0;
assign select_o[224] = (addr_i == 8'd224) ? 1 : 0;
assign select_o[225] = (addr_i == 8'd225) ? 1 : 0;
assign select_o[226] = (addr_i == 8'd226) ? 1 : 0;
assign select_o[227] = (addr_i == 8'd227) ? 1 : 0;
assign select_o[228] = (addr_i == 8'd228) ? 1 : 0;
assign select_o[229] = (addr_i == 8'd229) ? 1 : 0;
assign select_o[230] = (addr_i == 8'd230) ? 1 : 0;
assign select_o[231] = (addr_i == 8'd231) ? 1 : 0;
assign select_o[232] = (addr_i == 8'd232) ? 1 : 0;
assign select_o[233] = (addr_i == 8'd233) ? 1 : 0;
assign select_o[234] = (addr_i == 8'd234) ? 1 : 0;
assign select_o[235] = (addr_i == 8'd235) ? 1 : 0;
assign select_o[236] = (addr_i == 8'd236) ? 1 : 0;
assign select_o[237] = (addr_i == 8'd237) ? 1 : 0;
assign select_o[238] = (addr_i == 8'd238) ? 1 : 0;
assign select_o[239] = (addr_i == 8'd239) ? 1 : 0;
assign select_o[240] = (addr_i == 8'd240) ? 1 : 0;
assign select_o[241] = (addr_i == 8'd241) ? 1 : 0;
assign select_o[242] = (addr_i == 8'd242) ? 1 : 0;
assign select_o[243] = (addr_i == 8'd243) ? 1 : 0;
assign select_o[244] = (addr_i == 8'd244) ? 1 : 0;
assign select_o[245] = (addr_i == 8'd245) ? 1 : 0;
assign select_o[246] = (addr_i == 8'd246) ? 1 : 0;
assign select_o[247] = (addr_i == 8'd247) ? 1 : 0;
assign select_o[248] = (addr_i == 8'd248) ? 1 : 0;
assign select_o[249] = (addr_i == 8'd249) ? 1 : 0;
assign select_o[250] = (addr_i == 8'd250) ? 1 : 0;
assign select_o[251] = (addr_i == 8'd251) ? 1 : 0;
assign select_o[252] = (addr_i == 8'd252) ? 1 : 0;
assign select_o[253] = (addr_i == 8'd253) ? 1 : 0;
assign select_o[254] = (addr_i == 8'd254) ? 1 : 0;
assign select_o[255] = (addr_i == 8'd255) ? 1 : 0;
endmodule 