
module rbl(
	input  SLEEP,
	output CLK_RBL,
	output CLK_DIV,
	input  CLK
);

endmodule